magic
tech sky130A
magscale 1 2
timestamp 1669158044
<< obsli1 >>
rect 1104 2159 116840 161585
<< obsm1 >>
rect 290 892 117930 161616
<< metal2 >>
rect 478 163200 534 164000
rect 1398 163200 1454 164000
rect 2318 163200 2374 164000
rect 3238 163200 3294 164000
rect 4158 163200 4214 164000
rect 5078 163200 5134 164000
rect 5998 163200 6054 164000
rect 6918 163200 6974 164000
rect 7838 163200 7894 164000
rect 8758 163200 8814 164000
rect 9678 163200 9734 164000
rect 10598 163200 10654 164000
rect 11518 163200 11574 164000
rect 12438 163200 12494 164000
rect 13358 163200 13414 164000
rect 14278 163200 14334 164000
rect 15198 163200 15254 164000
rect 16118 163200 16174 164000
rect 17038 163200 17094 164000
rect 17958 163200 18014 164000
rect 18878 163200 18934 164000
rect 19798 163200 19854 164000
rect 20718 163200 20774 164000
rect 21638 163200 21694 164000
rect 22558 163200 22614 164000
rect 23478 163200 23534 164000
rect 24398 163200 24454 164000
rect 25318 163200 25374 164000
rect 26238 163200 26294 164000
rect 27158 163200 27214 164000
rect 28078 163200 28134 164000
rect 28998 163200 29054 164000
rect 29918 163200 29974 164000
rect 30838 163200 30894 164000
rect 31758 163200 31814 164000
rect 32678 163200 32734 164000
rect 33598 163200 33654 164000
rect 34518 163200 34574 164000
rect 35438 163200 35494 164000
rect 36358 163200 36414 164000
rect 37278 163200 37334 164000
rect 38198 163200 38254 164000
rect 39118 163200 39174 164000
rect 40038 163200 40094 164000
rect 40958 163200 41014 164000
rect 41878 163200 41934 164000
rect 42798 163200 42854 164000
rect 43718 163200 43774 164000
rect 44638 163200 44694 164000
rect 45558 163200 45614 164000
rect 46478 163200 46534 164000
rect 47398 163200 47454 164000
rect 48318 163200 48374 164000
rect 49238 163200 49294 164000
rect 50158 163200 50214 164000
rect 51078 163200 51134 164000
rect 51998 163200 52054 164000
rect 52918 163200 52974 164000
rect 53838 163200 53894 164000
rect 54758 163200 54814 164000
rect 55678 163200 55734 164000
rect 56598 163200 56654 164000
rect 57518 163200 57574 164000
rect 58438 163200 58494 164000
rect 59358 163200 59414 164000
rect 60278 163200 60334 164000
rect 61198 163200 61254 164000
rect 62118 163200 62174 164000
rect 63038 163200 63094 164000
rect 63958 163200 64014 164000
rect 64878 163200 64934 164000
rect 65798 163200 65854 164000
rect 66718 163200 66774 164000
rect 67638 163200 67694 164000
rect 68558 163200 68614 164000
rect 69478 163200 69534 164000
rect 70398 163200 70454 164000
rect 71318 163200 71374 164000
rect 72238 163200 72294 164000
rect 73158 163200 73214 164000
rect 74078 163200 74134 164000
rect 74998 163200 75054 164000
rect 75918 163200 75974 164000
rect 76838 163200 76894 164000
rect 77758 163200 77814 164000
rect 78678 163200 78734 164000
rect 79598 163200 79654 164000
rect 80518 163200 80574 164000
rect 81438 163200 81494 164000
rect 82358 163200 82414 164000
rect 83278 163200 83334 164000
rect 84198 163200 84254 164000
rect 85118 163200 85174 164000
rect 86038 163200 86094 164000
rect 86958 163200 87014 164000
rect 87878 163200 87934 164000
rect 88798 163200 88854 164000
rect 89718 163200 89774 164000
rect 90638 163200 90694 164000
rect 91558 163200 91614 164000
rect 92478 163200 92534 164000
rect 93398 163200 93454 164000
rect 94318 163200 94374 164000
rect 95238 163200 95294 164000
rect 96158 163200 96214 164000
rect 97078 163200 97134 164000
rect 97998 163200 98054 164000
rect 98918 163200 98974 164000
rect 99838 163200 99894 164000
rect 100758 163200 100814 164000
rect 101678 163200 101734 164000
rect 102598 163200 102654 164000
rect 103518 163200 103574 164000
rect 104438 163200 104494 164000
rect 105358 163200 105414 164000
rect 106278 163200 106334 164000
rect 107198 163200 107254 164000
rect 108118 163200 108174 164000
rect 109038 163200 109094 164000
rect 109958 163200 110014 164000
rect 110878 163200 110934 164000
rect 111798 163200 111854 164000
rect 112718 163200 112774 164000
rect 113638 163200 113694 164000
rect 114558 163200 114614 164000
rect 115478 163200 115534 164000
rect 116398 163200 116454 164000
rect 117318 163200 117374 164000
rect 294 0 350 800
rect 754 0 810 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17774 0 17830 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 20994 0 21050 800
rect 21454 0 21510 800
rect 21914 0 21970 800
rect 22374 0 22430 800
rect 22834 0 22890 800
rect 23294 0 23350 800
rect 23754 0 23810 800
rect 24214 0 24270 800
rect 24674 0 24730 800
rect 25134 0 25190 800
rect 25594 0 25650 800
rect 26054 0 26110 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27894 0 27950 800
rect 28354 0 28410 800
rect 28814 0 28870 800
rect 29274 0 29330 800
rect 29734 0 29790 800
rect 30194 0 30250 800
rect 30654 0 30710 800
rect 31114 0 31170 800
rect 31574 0 31630 800
rect 32034 0 32090 800
rect 32494 0 32550 800
rect 32954 0 33010 800
rect 33414 0 33470 800
rect 33874 0 33930 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36174 0 36230 800
rect 36634 0 36690 800
rect 37094 0 37150 800
rect 37554 0 37610 800
rect 38014 0 38070 800
rect 38474 0 38530 800
rect 38934 0 38990 800
rect 39394 0 39450 800
rect 39854 0 39910 800
rect 40314 0 40370 800
rect 40774 0 40830 800
rect 41234 0 41290 800
rect 41694 0 41750 800
rect 42154 0 42210 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 43994 0 44050 800
rect 44454 0 44510 800
rect 44914 0 44970 800
rect 45374 0 45430 800
rect 45834 0 45890 800
rect 46294 0 46350 800
rect 46754 0 46810 800
rect 47214 0 47270 800
rect 47674 0 47730 800
rect 48134 0 48190 800
rect 48594 0 48650 800
rect 49054 0 49110 800
rect 49514 0 49570 800
rect 49974 0 50030 800
rect 50434 0 50490 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53194 0 53250 800
rect 53654 0 53710 800
rect 54114 0 54170 800
rect 54574 0 54630 800
rect 55034 0 55090 800
rect 55494 0 55550 800
rect 55954 0 56010 800
rect 56414 0 56470 800
rect 56874 0 56930 800
rect 57334 0 57390 800
rect 57794 0 57850 800
rect 58254 0 58310 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
rect 60094 0 60150 800
rect 60554 0 60610 800
rect 61014 0 61070 800
rect 61474 0 61530 800
rect 61934 0 61990 800
rect 62394 0 62450 800
rect 62854 0 62910 800
rect 63314 0 63370 800
rect 63774 0 63830 800
rect 64234 0 64290 800
rect 64694 0 64750 800
rect 65154 0 65210 800
rect 65614 0 65670 800
rect 66074 0 66130 800
rect 66534 0 66590 800
rect 66994 0 67050 800
rect 67454 0 67510 800
rect 67914 0 67970 800
rect 68374 0 68430 800
rect 68834 0 68890 800
rect 69294 0 69350 800
rect 69754 0 69810 800
rect 70214 0 70270 800
rect 70674 0 70730 800
rect 71134 0 71190 800
rect 71594 0 71650 800
rect 72054 0 72110 800
rect 72514 0 72570 800
rect 72974 0 73030 800
rect 73434 0 73490 800
rect 73894 0 73950 800
rect 74354 0 74410 800
rect 74814 0 74870 800
rect 75274 0 75330 800
rect 75734 0 75790 800
rect 76194 0 76250 800
rect 76654 0 76710 800
rect 77114 0 77170 800
rect 77574 0 77630 800
rect 78034 0 78090 800
rect 78494 0 78550 800
rect 78954 0 79010 800
rect 79414 0 79470 800
rect 79874 0 79930 800
rect 80334 0 80390 800
rect 80794 0 80850 800
rect 81254 0 81310 800
rect 81714 0 81770 800
rect 82174 0 82230 800
rect 82634 0 82690 800
rect 83094 0 83150 800
rect 83554 0 83610 800
rect 84014 0 84070 800
rect 84474 0 84530 800
rect 84934 0 84990 800
rect 85394 0 85450 800
rect 85854 0 85910 800
rect 86314 0 86370 800
rect 86774 0 86830 800
rect 87234 0 87290 800
rect 87694 0 87750 800
rect 88154 0 88210 800
rect 88614 0 88670 800
rect 89074 0 89130 800
rect 89534 0 89590 800
rect 89994 0 90050 800
rect 90454 0 90510 800
rect 90914 0 90970 800
rect 91374 0 91430 800
rect 91834 0 91890 800
rect 92294 0 92350 800
rect 92754 0 92810 800
rect 93214 0 93270 800
rect 93674 0 93730 800
rect 94134 0 94190 800
rect 94594 0 94650 800
rect 95054 0 95110 800
rect 95514 0 95570 800
rect 95974 0 96030 800
rect 96434 0 96490 800
rect 96894 0 96950 800
rect 97354 0 97410 800
rect 97814 0 97870 800
rect 98274 0 98330 800
rect 98734 0 98790 800
rect 99194 0 99250 800
rect 99654 0 99710 800
rect 100114 0 100170 800
rect 100574 0 100630 800
rect 101034 0 101090 800
rect 101494 0 101550 800
rect 101954 0 102010 800
rect 102414 0 102470 800
rect 102874 0 102930 800
rect 103334 0 103390 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104714 0 104770 800
rect 105174 0 105230 800
rect 105634 0 105690 800
rect 106094 0 106150 800
rect 106554 0 106610 800
rect 107014 0 107070 800
rect 107474 0 107530 800
rect 107934 0 107990 800
rect 108394 0 108450 800
rect 108854 0 108910 800
rect 109314 0 109370 800
rect 109774 0 109830 800
rect 110234 0 110290 800
rect 110694 0 110750 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 112074 0 112130 800
rect 112534 0 112590 800
rect 112994 0 113050 800
rect 113454 0 113510 800
rect 113914 0 113970 800
rect 114374 0 114430 800
rect 114834 0 114890 800
rect 115294 0 115350 800
rect 115754 0 115810 800
rect 116214 0 116270 800
rect 116674 0 116730 800
rect 117134 0 117190 800
rect 117594 0 117650 800
<< obsm2 >>
rect 296 163144 422 163282
rect 590 163144 1342 163282
rect 1510 163144 2262 163282
rect 2430 163144 3182 163282
rect 3350 163144 4102 163282
rect 4270 163144 5022 163282
rect 5190 163144 5942 163282
rect 6110 163144 6862 163282
rect 7030 163144 7782 163282
rect 7950 163144 8702 163282
rect 8870 163144 9622 163282
rect 9790 163144 10542 163282
rect 10710 163144 11462 163282
rect 11630 163144 12382 163282
rect 12550 163144 13302 163282
rect 13470 163144 14222 163282
rect 14390 163144 15142 163282
rect 15310 163144 16062 163282
rect 16230 163144 16982 163282
rect 17150 163144 17902 163282
rect 18070 163144 18822 163282
rect 18990 163144 19742 163282
rect 19910 163144 20662 163282
rect 20830 163144 21582 163282
rect 21750 163144 22502 163282
rect 22670 163144 23422 163282
rect 23590 163144 24342 163282
rect 24510 163144 25262 163282
rect 25430 163144 26182 163282
rect 26350 163144 27102 163282
rect 27270 163144 28022 163282
rect 28190 163144 28942 163282
rect 29110 163144 29862 163282
rect 30030 163144 30782 163282
rect 30950 163144 31702 163282
rect 31870 163144 32622 163282
rect 32790 163144 33542 163282
rect 33710 163144 34462 163282
rect 34630 163144 35382 163282
rect 35550 163144 36302 163282
rect 36470 163144 37222 163282
rect 37390 163144 38142 163282
rect 38310 163144 39062 163282
rect 39230 163144 39982 163282
rect 40150 163144 40902 163282
rect 41070 163144 41822 163282
rect 41990 163144 42742 163282
rect 42910 163144 43662 163282
rect 43830 163144 44582 163282
rect 44750 163144 45502 163282
rect 45670 163144 46422 163282
rect 46590 163144 47342 163282
rect 47510 163144 48262 163282
rect 48430 163144 49182 163282
rect 49350 163144 50102 163282
rect 50270 163144 51022 163282
rect 51190 163144 51942 163282
rect 52110 163144 52862 163282
rect 53030 163144 53782 163282
rect 53950 163144 54702 163282
rect 54870 163144 55622 163282
rect 55790 163144 56542 163282
rect 56710 163144 57462 163282
rect 57630 163144 58382 163282
rect 58550 163144 59302 163282
rect 59470 163144 60222 163282
rect 60390 163144 61142 163282
rect 61310 163144 62062 163282
rect 62230 163144 62982 163282
rect 63150 163144 63902 163282
rect 64070 163144 64822 163282
rect 64990 163144 65742 163282
rect 65910 163144 66662 163282
rect 66830 163144 67582 163282
rect 67750 163144 68502 163282
rect 68670 163144 69422 163282
rect 69590 163144 70342 163282
rect 70510 163144 71262 163282
rect 71430 163144 72182 163282
rect 72350 163144 73102 163282
rect 73270 163144 74022 163282
rect 74190 163144 74942 163282
rect 75110 163144 75862 163282
rect 76030 163144 76782 163282
rect 76950 163144 77702 163282
rect 77870 163144 78622 163282
rect 78790 163144 79542 163282
rect 79710 163144 80462 163282
rect 80630 163144 81382 163282
rect 81550 163144 82302 163282
rect 82470 163144 83222 163282
rect 83390 163144 84142 163282
rect 84310 163144 85062 163282
rect 85230 163144 85982 163282
rect 86150 163144 86902 163282
rect 87070 163144 87822 163282
rect 87990 163144 88742 163282
rect 88910 163144 89662 163282
rect 89830 163144 90582 163282
rect 90750 163144 91502 163282
rect 91670 163144 92422 163282
rect 92590 163144 93342 163282
rect 93510 163144 94262 163282
rect 94430 163144 95182 163282
rect 95350 163144 96102 163282
rect 96270 163144 97022 163282
rect 97190 163144 97942 163282
rect 98110 163144 98862 163282
rect 99030 163144 99782 163282
rect 99950 163144 100702 163282
rect 100870 163144 101622 163282
rect 101790 163144 102542 163282
rect 102710 163144 103462 163282
rect 103630 163144 104382 163282
rect 104550 163144 105302 163282
rect 105470 163144 106222 163282
rect 106390 163144 107142 163282
rect 107310 163144 108062 163282
rect 108230 163144 108982 163282
rect 109150 163144 109902 163282
rect 110070 163144 110822 163282
rect 110990 163144 111742 163282
rect 111910 163144 112662 163282
rect 112830 163144 113582 163282
rect 113750 163144 114502 163282
rect 114670 163144 115422 163282
rect 115590 163144 116342 163282
rect 116510 163144 117262 163282
rect 117430 163144 117924 163282
rect 296 856 117924 163144
rect 406 734 698 856
rect 866 734 1158 856
rect 1326 734 1618 856
rect 1786 734 2078 856
rect 2246 734 2538 856
rect 2706 734 2998 856
rect 3166 734 3458 856
rect 3626 734 3918 856
rect 4086 734 4378 856
rect 4546 734 4838 856
rect 5006 734 5298 856
rect 5466 734 5758 856
rect 5926 734 6218 856
rect 6386 734 6678 856
rect 6846 734 7138 856
rect 7306 734 7598 856
rect 7766 734 8058 856
rect 8226 734 8518 856
rect 8686 734 8978 856
rect 9146 734 9438 856
rect 9606 734 9898 856
rect 10066 734 10358 856
rect 10526 734 10818 856
rect 10986 734 11278 856
rect 11446 734 11738 856
rect 11906 734 12198 856
rect 12366 734 12658 856
rect 12826 734 13118 856
rect 13286 734 13578 856
rect 13746 734 14038 856
rect 14206 734 14498 856
rect 14666 734 14958 856
rect 15126 734 15418 856
rect 15586 734 15878 856
rect 16046 734 16338 856
rect 16506 734 16798 856
rect 16966 734 17258 856
rect 17426 734 17718 856
rect 17886 734 18178 856
rect 18346 734 18638 856
rect 18806 734 19098 856
rect 19266 734 19558 856
rect 19726 734 20018 856
rect 20186 734 20478 856
rect 20646 734 20938 856
rect 21106 734 21398 856
rect 21566 734 21858 856
rect 22026 734 22318 856
rect 22486 734 22778 856
rect 22946 734 23238 856
rect 23406 734 23698 856
rect 23866 734 24158 856
rect 24326 734 24618 856
rect 24786 734 25078 856
rect 25246 734 25538 856
rect 25706 734 25998 856
rect 26166 734 26458 856
rect 26626 734 26918 856
rect 27086 734 27378 856
rect 27546 734 27838 856
rect 28006 734 28298 856
rect 28466 734 28758 856
rect 28926 734 29218 856
rect 29386 734 29678 856
rect 29846 734 30138 856
rect 30306 734 30598 856
rect 30766 734 31058 856
rect 31226 734 31518 856
rect 31686 734 31978 856
rect 32146 734 32438 856
rect 32606 734 32898 856
rect 33066 734 33358 856
rect 33526 734 33818 856
rect 33986 734 34278 856
rect 34446 734 34738 856
rect 34906 734 35198 856
rect 35366 734 35658 856
rect 35826 734 36118 856
rect 36286 734 36578 856
rect 36746 734 37038 856
rect 37206 734 37498 856
rect 37666 734 37958 856
rect 38126 734 38418 856
rect 38586 734 38878 856
rect 39046 734 39338 856
rect 39506 734 39798 856
rect 39966 734 40258 856
rect 40426 734 40718 856
rect 40886 734 41178 856
rect 41346 734 41638 856
rect 41806 734 42098 856
rect 42266 734 42558 856
rect 42726 734 43018 856
rect 43186 734 43478 856
rect 43646 734 43938 856
rect 44106 734 44398 856
rect 44566 734 44858 856
rect 45026 734 45318 856
rect 45486 734 45778 856
rect 45946 734 46238 856
rect 46406 734 46698 856
rect 46866 734 47158 856
rect 47326 734 47618 856
rect 47786 734 48078 856
rect 48246 734 48538 856
rect 48706 734 48998 856
rect 49166 734 49458 856
rect 49626 734 49918 856
rect 50086 734 50378 856
rect 50546 734 50838 856
rect 51006 734 51298 856
rect 51466 734 51758 856
rect 51926 734 52218 856
rect 52386 734 52678 856
rect 52846 734 53138 856
rect 53306 734 53598 856
rect 53766 734 54058 856
rect 54226 734 54518 856
rect 54686 734 54978 856
rect 55146 734 55438 856
rect 55606 734 55898 856
rect 56066 734 56358 856
rect 56526 734 56818 856
rect 56986 734 57278 856
rect 57446 734 57738 856
rect 57906 734 58198 856
rect 58366 734 58658 856
rect 58826 734 59118 856
rect 59286 734 59578 856
rect 59746 734 60038 856
rect 60206 734 60498 856
rect 60666 734 60958 856
rect 61126 734 61418 856
rect 61586 734 61878 856
rect 62046 734 62338 856
rect 62506 734 62798 856
rect 62966 734 63258 856
rect 63426 734 63718 856
rect 63886 734 64178 856
rect 64346 734 64638 856
rect 64806 734 65098 856
rect 65266 734 65558 856
rect 65726 734 66018 856
rect 66186 734 66478 856
rect 66646 734 66938 856
rect 67106 734 67398 856
rect 67566 734 67858 856
rect 68026 734 68318 856
rect 68486 734 68778 856
rect 68946 734 69238 856
rect 69406 734 69698 856
rect 69866 734 70158 856
rect 70326 734 70618 856
rect 70786 734 71078 856
rect 71246 734 71538 856
rect 71706 734 71998 856
rect 72166 734 72458 856
rect 72626 734 72918 856
rect 73086 734 73378 856
rect 73546 734 73838 856
rect 74006 734 74298 856
rect 74466 734 74758 856
rect 74926 734 75218 856
rect 75386 734 75678 856
rect 75846 734 76138 856
rect 76306 734 76598 856
rect 76766 734 77058 856
rect 77226 734 77518 856
rect 77686 734 77978 856
rect 78146 734 78438 856
rect 78606 734 78898 856
rect 79066 734 79358 856
rect 79526 734 79818 856
rect 79986 734 80278 856
rect 80446 734 80738 856
rect 80906 734 81198 856
rect 81366 734 81658 856
rect 81826 734 82118 856
rect 82286 734 82578 856
rect 82746 734 83038 856
rect 83206 734 83498 856
rect 83666 734 83958 856
rect 84126 734 84418 856
rect 84586 734 84878 856
rect 85046 734 85338 856
rect 85506 734 85798 856
rect 85966 734 86258 856
rect 86426 734 86718 856
rect 86886 734 87178 856
rect 87346 734 87638 856
rect 87806 734 88098 856
rect 88266 734 88558 856
rect 88726 734 89018 856
rect 89186 734 89478 856
rect 89646 734 89938 856
rect 90106 734 90398 856
rect 90566 734 90858 856
rect 91026 734 91318 856
rect 91486 734 91778 856
rect 91946 734 92238 856
rect 92406 734 92698 856
rect 92866 734 93158 856
rect 93326 734 93618 856
rect 93786 734 94078 856
rect 94246 734 94538 856
rect 94706 734 94998 856
rect 95166 734 95458 856
rect 95626 734 95918 856
rect 96086 734 96378 856
rect 96546 734 96838 856
rect 97006 734 97298 856
rect 97466 734 97758 856
rect 97926 734 98218 856
rect 98386 734 98678 856
rect 98846 734 99138 856
rect 99306 734 99598 856
rect 99766 734 100058 856
rect 100226 734 100518 856
rect 100686 734 100978 856
rect 101146 734 101438 856
rect 101606 734 101898 856
rect 102066 734 102358 856
rect 102526 734 102818 856
rect 102986 734 103278 856
rect 103446 734 103738 856
rect 103906 734 104198 856
rect 104366 734 104658 856
rect 104826 734 105118 856
rect 105286 734 105578 856
rect 105746 734 106038 856
rect 106206 734 106498 856
rect 106666 734 106958 856
rect 107126 734 107418 856
rect 107586 734 107878 856
rect 108046 734 108338 856
rect 108506 734 108798 856
rect 108966 734 109258 856
rect 109426 734 109718 856
rect 109886 734 110178 856
rect 110346 734 110638 856
rect 110806 734 111098 856
rect 111266 734 111558 856
rect 111726 734 112018 856
rect 112186 734 112478 856
rect 112646 734 112938 856
rect 113106 734 113398 856
rect 113566 734 113858 856
rect 114026 734 114318 856
rect 114486 734 114778 856
rect 114946 734 115238 856
rect 115406 734 115698 856
rect 115866 734 116158 856
rect 116326 734 116618 856
rect 116786 734 117078 856
rect 117246 734 117538 856
rect 117706 734 117924 856
<< metal3 >>
rect 117200 161848 118000 161968
rect 0 159944 800 160064
rect 117200 158448 118000 158568
rect 117200 155048 118000 155168
rect 0 154368 800 154488
rect 117200 151648 118000 151768
rect 0 148792 800 148912
rect 117200 148248 118000 148368
rect 117200 144848 118000 144968
rect 0 143216 800 143336
rect 117200 141448 118000 141568
rect 117200 138048 118000 138168
rect 0 137640 800 137760
rect 117200 134648 118000 134768
rect 0 132064 800 132184
rect 117200 131248 118000 131368
rect 117200 127848 118000 127968
rect 0 126488 800 126608
rect 117200 124448 118000 124568
rect 0 120912 800 121032
rect 117200 121048 118000 121168
rect 117200 117648 118000 117768
rect 0 115336 800 115456
rect 117200 114248 118000 114368
rect 117200 110848 118000 110968
rect 0 109760 800 109880
rect 117200 107448 118000 107568
rect 0 104184 800 104304
rect 117200 104048 118000 104168
rect 117200 100648 118000 100768
rect 0 98608 800 98728
rect 117200 97248 118000 97368
rect 117200 93848 118000 93968
rect 0 93032 800 93152
rect 117200 90448 118000 90568
rect 0 87456 800 87576
rect 117200 87048 118000 87168
rect 117200 83648 118000 83768
rect 0 81880 800 82000
rect 117200 80248 118000 80368
rect 117200 76848 118000 76968
rect 0 76304 800 76424
rect 117200 73448 118000 73568
rect 0 70728 800 70848
rect 117200 70048 118000 70168
rect 117200 66648 118000 66768
rect 0 65152 800 65272
rect 117200 63248 118000 63368
rect 117200 59848 118000 59968
rect 0 59576 800 59696
rect 117200 56448 118000 56568
rect 0 54000 800 54120
rect 117200 53048 118000 53168
rect 117200 49648 118000 49768
rect 0 48424 800 48544
rect 117200 46248 118000 46368
rect 0 42848 800 42968
rect 117200 42848 118000 42968
rect 117200 39448 118000 39568
rect 0 37272 800 37392
rect 117200 36048 118000 36168
rect 117200 32648 118000 32768
rect 0 31696 800 31816
rect 117200 29248 118000 29368
rect 0 26120 800 26240
rect 117200 25848 118000 25968
rect 117200 22448 118000 22568
rect 0 20544 800 20664
rect 117200 19048 118000 19168
rect 117200 15648 118000 15768
rect 0 14968 800 15088
rect 117200 12248 118000 12368
rect 0 9392 800 9512
rect 117200 8848 118000 8968
rect 117200 5448 118000 5568
rect 0 3816 800 3936
rect 117200 2048 118000 2168
<< obsm3 >>
rect 800 161768 117120 161940
rect 800 160144 117200 161768
rect 880 159864 117200 160144
rect 800 158648 117200 159864
rect 800 158368 117120 158648
rect 800 155248 117200 158368
rect 800 154968 117120 155248
rect 800 154568 117200 154968
rect 880 154288 117200 154568
rect 800 151848 117200 154288
rect 800 151568 117120 151848
rect 800 148992 117200 151568
rect 880 148712 117200 148992
rect 800 148448 117200 148712
rect 800 148168 117120 148448
rect 800 145048 117200 148168
rect 800 144768 117120 145048
rect 800 143416 117200 144768
rect 880 143136 117200 143416
rect 800 141648 117200 143136
rect 800 141368 117120 141648
rect 800 138248 117200 141368
rect 800 137968 117120 138248
rect 800 137840 117200 137968
rect 880 137560 117200 137840
rect 800 134848 117200 137560
rect 800 134568 117120 134848
rect 800 132264 117200 134568
rect 880 131984 117200 132264
rect 800 131448 117200 131984
rect 800 131168 117120 131448
rect 800 128048 117200 131168
rect 800 127768 117120 128048
rect 800 126688 117200 127768
rect 880 126408 117200 126688
rect 800 124648 117200 126408
rect 800 124368 117120 124648
rect 800 121248 117200 124368
rect 800 121112 117120 121248
rect 880 120968 117120 121112
rect 880 120832 117200 120968
rect 800 117848 117200 120832
rect 800 117568 117120 117848
rect 800 115536 117200 117568
rect 880 115256 117200 115536
rect 800 114448 117200 115256
rect 800 114168 117120 114448
rect 800 111048 117200 114168
rect 800 110768 117120 111048
rect 800 109960 117200 110768
rect 880 109680 117200 109960
rect 800 107648 117200 109680
rect 800 107368 117120 107648
rect 800 104384 117200 107368
rect 880 104248 117200 104384
rect 880 104104 117120 104248
rect 800 103968 117120 104104
rect 800 100848 117200 103968
rect 800 100568 117120 100848
rect 800 98808 117200 100568
rect 880 98528 117200 98808
rect 800 97448 117200 98528
rect 800 97168 117120 97448
rect 800 94048 117200 97168
rect 800 93768 117120 94048
rect 800 93232 117200 93768
rect 880 92952 117200 93232
rect 800 90648 117200 92952
rect 800 90368 117120 90648
rect 800 87656 117200 90368
rect 880 87376 117200 87656
rect 800 87248 117200 87376
rect 800 86968 117120 87248
rect 800 83848 117200 86968
rect 800 83568 117120 83848
rect 800 82080 117200 83568
rect 880 81800 117200 82080
rect 800 80448 117200 81800
rect 800 80168 117120 80448
rect 800 77048 117200 80168
rect 800 76768 117120 77048
rect 800 76504 117200 76768
rect 880 76224 117200 76504
rect 800 73648 117200 76224
rect 800 73368 117120 73648
rect 800 70928 117200 73368
rect 880 70648 117200 70928
rect 800 70248 117200 70648
rect 800 69968 117120 70248
rect 800 66848 117200 69968
rect 800 66568 117120 66848
rect 800 65352 117200 66568
rect 880 65072 117200 65352
rect 800 63448 117200 65072
rect 800 63168 117120 63448
rect 800 60048 117200 63168
rect 800 59776 117120 60048
rect 880 59768 117120 59776
rect 880 59496 117200 59768
rect 800 56648 117200 59496
rect 800 56368 117120 56648
rect 800 54200 117200 56368
rect 880 53920 117200 54200
rect 800 53248 117200 53920
rect 800 52968 117120 53248
rect 800 49848 117200 52968
rect 800 49568 117120 49848
rect 800 48624 117200 49568
rect 880 48344 117200 48624
rect 800 46448 117200 48344
rect 800 46168 117120 46448
rect 800 43048 117200 46168
rect 880 42768 117120 43048
rect 800 39648 117200 42768
rect 800 39368 117120 39648
rect 800 37472 117200 39368
rect 880 37192 117200 37472
rect 800 36248 117200 37192
rect 800 35968 117120 36248
rect 800 32848 117200 35968
rect 800 32568 117120 32848
rect 800 31896 117200 32568
rect 880 31616 117200 31896
rect 800 29448 117200 31616
rect 800 29168 117120 29448
rect 800 26320 117200 29168
rect 880 26048 117200 26320
rect 880 26040 117120 26048
rect 800 25768 117120 26040
rect 800 22648 117200 25768
rect 800 22368 117120 22648
rect 800 20744 117200 22368
rect 880 20464 117200 20744
rect 800 19248 117200 20464
rect 800 18968 117120 19248
rect 800 15848 117200 18968
rect 800 15568 117120 15848
rect 800 15168 117200 15568
rect 880 14888 117200 15168
rect 800 12448 117200 14888
rect 800 12168 117120 12448
rect 800 9592 117200 12168
rect 880 9312 117200 9592
rect 800 9048 117200 9312
rect 800 8768 117120 9048
rect 800 5648 117200 8768
rect 800 5368 117120 5648
rect 800 4016 117200 5368
rect 880 3736 117200 4016
rect 800 2248 117200 3736
rect 800 1968 117120 2248
rect 800 1803 117200 1968
<< metal4 >>
rect 4208 2128 4528 161616
rect 19568 2128 19888 161616
rect 34928 2128 35248 161616
rect 50288 2128 50608 161616
rect 65648 2128 65968 161616
rect 81008 2128 81328 161616
rect 96368 2128 96688 161616
rect 111728 2128 112048 161616
<< obsm4 >>
rect 1899 161696 116045 161941
rect 1899 2048 4128 161696
rect 4608 2048 19488 161696
rect 19968 2048 34848 161696
rect 35328 2048 50208 161696
rect 50688 2048 65568 161696
rect 66048 2048 80928 161696
rect 81408 2048 96288 161696
rect 96768 2048 111648 161696
rect 112128 2048 116045 161696
rect 1899 1803 116045 2048
<< labels >>
rlabel metal3 s 0 159944 800 160064 6 clk
port 1 nsew signal input
rlabel metal3 s 117200 2048 118000 2168 6 raddr0[0]
port 2 nsew signal input
rlabel metal3 s 117200 29248 118000 29368 6 raddr0[1]
port 3 nsew signal input
rlabel metal3 s 117200 56448 118000 56568 6 raddr0[2]
port 4 nsew signal input
rlabel metal3 s 117200 83648 118000 83768 6 raddr0[3]
port 5 nsew signal input
rlabel metal3 s 117200 110848 118000 110968 6 raddr0[4]
port 6 nsew signal input
rlabel metal3 s 117200 138048 118000 138168 6 raddr0[5]
port 7 nsew signal input
rlabel metal3 s 117200 5448 118000 5568 6 raddr1[0]
port 8 nsew signal input
rlabel metal3 s 117200 32648 118000 32768 6 raddr1[1]
port 9 nsew signal input
rlabel metal3 s 117200 59848 118000 59968 6 raddr1[2]
port 10 nsew signal input
rlabel metal3 s 117200 87048 118000 87168 6 raddr1[3]
port 11 nsew signal input
rlabel metal3 s 117200 114248 118000 114368 6 raddr1[4]
port 12 nsew signal input
rlabel metal3 s 117200 141448 118000 141568 6 raddr1[5]
port 13 nsew signal input
rlabel metal3 s 117200 8848 118000 8968 6 raddr2[0]
port 14 nsew signal input
rlabel metal3 s 117200 36048 118000 36168 6 raddr2[1]
port 15 nsew signal input
rlabel metal3 s 117200 63248 118000 63368 6 raddr2[2]
port 16 nsew signal input
rlabel metal3 s 117200 90448 118000 90568 6 raddr2[3]
port 17 nsew signal input
rlabel metal3 s 117200 117648 118000 117768 6 raddr2[4]
port 18 nsew signal input
rlabel metal3 s 117200 144848 118000 144968 6 raddr2[5]
port 19 nsew signal input
rlabel metal3 s 117200 12248 118000 12368 6 raddr3[0]
port 20 nsew signal input
rlabel metal3 s 117200 39448 118000 39568 6 raddr3[1]
port 21 nsew signal input
rlabel metal3 s 117200 66648 118000 66768 6 raddr3[2]
port 22 nsew signal input
rlabel metal3 s 117200 93848 118000 93968 6 raddr3[3]
port 23 nsew signal input
rlabel metal3 s 117200 121048 118000 121168 6 raddr3[4]
port 24 nsew signal input
rlabel metal3 s 117200 148248 118000 148368 6 raddr3[5]
port 25 nsew signal input
rlabel metal3 s 117200 15648 118000 15768 6 raddr4[0]
port 26 nsew signal input
rlabel metal3 s 117200 42848 118000 42968 6 raddr4[1]
port 27 nsew signal input
rlabel metal3 s 117200 70048 118000 70168 6 raddr4[2]
port 28 nsew signal input
rlabel metal3 s 117200 97248 118000 97368 6 raddr4[3]
port 29 nsew signal input
rlabel metal3 s 117200 124448 118000 124568 6 raddr4[4]
port 30 nsew signal input
rlabel metal3 s 117200 151648 118000 151768 6 raddr4[5]
port 31 nsew signal input
rlabel metal3 s 117200 19048 118000 19168 6 raddr5[0]
port 32 nsew signal input
rlabel metal3 s 117200 46248 118000 46368 6 raddr5[1]
port 33 nsew signal input
rlabel metal3 s 117200 73448 118000 73568 6 raddr5[2]
port 34 nsew signal input
rlabel metal3 s 117200 100648 118000 100768 6 raddr5[3]
port 35 nsew signal input
rlabel metal3 s 117200 127848 118000 127968 6 raddr5[4]
port 36 nsew signal input
rlabel metal3 s 117200 155048 118000 155168 6 raddr5[5]
port 37 nsew signal input
rlabel metal3 s 117200 22448 118000 22568 6 raddr6[0]
port 38 nsew signal input
rlabel metal3 s 117200 49648 118000 49768 6 raddr6[1]
port 39 nsew signal input
rlabel metal3 s 117200 76848 118000 76968 6 raddr6[2]
port 40 nsew signal input
rlabel metal3 s 117200 104048 118000 104168 6 raddr6[3]
port 41 nsew signal input
rlabel metal3 s 117200 131248 118000 131368 6 raddr6[4]
port 42 nsew signal input
rlabel metal3 s 117200 158448 118000 158568 6 raddr6[5]
port 43 nsew signal input
rlabel metal3 s 117200 25848 118000 25968 6 raddr7[0]
port 44 nsew signal input
rlabel metal3 s 117200 53048 118000 53168 6 raddr7[1]
port 45 nsew signal input
rlabel metal3 s 117200 80248 118000 80368 6 raddr7[2]
port 46 nsew signal input
rlabel metal3 s 117200 107448 118000 107568 6 raddr7[3]
port 47 nsew signal input
rlabel metal3 s 117200 134648 118000 134768 6 raddr7[4]
port 48 nsew signal input
rlabel metal3 s 117200 161848 118000 161968 6 raddr7[5]
port 49 nsew signal input
rlabel metal2 s 294 0 350 800 6 rdata0[0]
port 50 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 rdata0[10]
port 51 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 rdata0[11]
port 52 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 rdata0[12]
port 53 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 rdata0[13]
port 54 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 rdata0[14]
port 55 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 rdata0[15]
port 56 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 rdata0[16]
port 57 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 rdata0[17]
port 58 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 rdata0[18]
port 59 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 rdata0[19]
port 60 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 rdata0[1]
port 61 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 rdata0[20]
port 62 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 rdata0[21]
port 63 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 rdata0[22]
port 64 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 rdata0[23]
port 65 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 rdata0[24]
port 66 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 rdata0[25]
port 67 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 rdata0[26]
port 68 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 rdata0[27]
port 69 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 rdata0[28]
port 70 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 rdata0[29]
port 71 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 rdata0[2]
port 72 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 rdata0[30]
port 73 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 rdata0[31]
port 74 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 rdata0[3]
port 75 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 rdata0[4]
port 76 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 rdata0[5]
port 77 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 rdata0[6]
port 78 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 rdata0[7]
port 79 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 rdata0[8]
port 80 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 rdata0[9]
port 81 nsew signal output
rlabel metal2 s 754 0 810 800 6 rdata1[0]
port 82 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 rdata1[10]
port 83 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 rdata1[11]
port 84 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 rdata1[12]
port 85 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 rdata1[13]
port 86 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 rdata1[14]
port 87 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 rdata1[15]
port 88 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 rdata1[16]
port 89 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 rdata1[17]
port 90 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 rdata1[18]
port 91 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 rdata1[19]
port 92 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 rdata1[1]
port 93 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 rdata1[20]
port 94 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 rdata1[21]
port 95 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 rdata1[22]
port 96 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 rdata1[23]
port 97 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 rdata1[24]
port 98 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 rdata1[25]
port 99 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 rdata1[26]
port 100 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 rdata1[27]
port 101 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 rdata1[28]
port 102 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 rdata1[29]
port 103 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 rdata1[2]
port 104 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 rdata1[30]
port 105 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 rdata1[31]
port 106 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 rdata1[3]
port 107 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 rdata1[4]
port 108 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 rdata1[5]
port 109 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 rdata1[6]
port 110 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 rdata1[7]
port 111 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 rdata1[8]
port 112 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 rdata1[9]
port 113 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 rdata2[0]
port 114 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 rdata2[10]
port 115 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 rdata2[11]
port 116 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 rdata2[12]
port 117 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 rdata2[13]
port 118 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 rdata2[14]
port 119 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 rdata2[15]
port 120 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 rdata2[16]
port 121 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 rdata2[17]
port 122 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 rdata2[18]
port 123 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 rdata2[19]
port 124 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 rdata2[1]
port 125 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 rdata2[20]
port 126 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 rdata2[21]
port 127 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 rdata2[22]
port 128 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 rdata2[23]
port 129 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 rdata2[24]
port 130 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 rdata2[25]
port 131 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 rdata2[26]
port 132 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 rdata2[27]
port 133 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 rdata2[28]
port 134 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 rdata2[29]
port 135 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 rdata2[2]
port 136 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 rdata2[30]
port 137 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 rdata2[31]
port 138 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 rdata2[3]
port 139 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 rdata2[4]
port 140 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 rdata2[5]
port 141 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 rdata2[6]
port 142 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 rdata2[7]
port 143 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 rdata2[8]
port 144 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 rdata2[9]
port 145 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 rdata3[0]
port 146 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 rdata3[10]
port 147 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 rdata3[11]
port 148 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 rdata3[12]
port 149 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 rdata3[13]
port 150 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 rdata3[14]
port 151 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 rdata3[15]
port 152 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 rdata3[16]
port 153 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 rdata3[17]
port 154 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 rdata3[18]
port 155 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 rdata3[19]
port 156 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 rdata3[1]
port 157 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 rdata3[20]
port 158 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 rdata3[21]
port 159 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 rdata3[22]
port 160 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 rdata3[23]
port 161 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 rdata3[24]
port 162 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 rdata3[25]
port 163 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 rdata3[26]
port 164 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 rdata3[27]
port 165 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 rdata3[28]
port 166 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 rdata3[29]
port 167 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 rdata3[2]
port 168 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 rdata3[30]
port 169 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 rdata3[31]
port 170 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 rdata3[3]
port 171 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 rdata3[4]
port 172 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 rdata3[5]
port 173 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 rdata3[6]
port 174 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 rdata3[7]
port 175 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 rdata3[8]
port 176 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 rdata3[9]
port 177 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 rdata4[0]
port 178 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 rdata4[10]
port 179 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 rdata4[11]
port 180 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 rdata4[12]
port 181 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 rdata4[13]
port 182 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 rdata4[14]
port 183 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 rdata4[15]
port 184 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 rdata4[16]
port 185 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 rdata4[17]
port 186 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 rdata4[18]
port 187 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 rdata4[19]
port 188 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 rdata4[1]
port 189 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 rdata4[20]
port 190 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 rdata4[21]
port 191 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 rdata4[22]
port 192 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 rdata4[23]
port 193 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 rdata4[24]
port 194 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 rdata4[25]
port 195 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 rdata4[26]
port 196 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 rdata4[27]
port 197 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 rdata4[28]
port 198 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 rdata4[29]
port 199 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 rdata4[2]
port 200 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 rdata4[30]
port 201 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 rdata4[31]
port 202 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 rdata4[3]
port 203 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 rdata4[4]
port 204 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 rdata4[5]
port 205 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 rdata4[6]
port 206 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 rdata4[7]
port 207 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 rdata4[8]
port 208 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 rdata4[9]
port 209 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 rdata5[0]
port 210 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 rdata5[10]
port 211 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 rdata5[11]
port 212 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 rdata5[12]
port 213 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 rdata5[13]
port 214 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 rdata5[14]
port 215 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 rdata5[15]
port 216 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 rdata5[16]
port 217 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 rdata5[17]
port 218 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 rdata5[18]
port 219 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 rdata5[19]
port 220 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 rdata5[1]
port 221 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 rdata5[20]
port 222 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 rdata5[21]
port 223 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 rdata5[22]
port 224 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 rdata5[23]
port 225 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 rdata5[24]
port 226 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 rdata5[25]
port 227 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 rdata5[26]
port 228 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 rdata5[27]
port 229 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 rdata5[28]
port 230 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 rdata5[29]
port 231 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 rdata5[2]
port 232 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 rdata5[30]
port 233 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 rdata5[31]
port 234 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 rdata5[3]
port 235 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 rdata5[4]
port 236 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 rdata5[5]
port 237 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 rdata5[6]
port 238 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 rdata5[7]
port 239 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 rdata5[8]
port 240 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 rdata5[9]
port 241 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 rdata6[0]
port 242 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 rdata6[10]
port 243 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 rdata6[11]
port 244 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 rdata6[12]
port 245 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 rdata6[13]
port 246 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 rdata6[14]
port 247 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 rdata6[15]
port 248 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 rdata6[16]
port 249 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 rdata6[17]
port 250 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 rdata6[18]
port 251 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 rdata6[19]
port 252 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 rdata6[1]
port 253 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 rdata6[20]
port 254 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 rdata6[21]
port 255 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 rdata6[22]
port 256 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 rdata6[23]
port 257 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 rdata6[24]
port 258 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 rdata6[25]
port 259 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 rdata6[26]
port 260 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 rdata6[27]
port 261 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 rdata6[28]
port 262 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 rdata6[29]
port 263 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 rdata6[2]
port 264 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 rdata6[30]
port 265 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 rdata6[31]
port 266 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 rdata6[3]
port 267 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 rdata6[4]
port 268 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 rdata6[5]
port 269 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 rdata6[6]
port 270 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 rdata6[7]
port 271 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 rdata6[8]
port 272 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 rdata6[9]
port 273 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 rdata7[0]
port 274 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 rdata7[10]
port 275 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 rdata7[11]
port 276 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 rdata7[12]
port 277 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 rdata7[13]
port 278 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 rdata7[14]
port 279 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 rdata7[15]
port 280 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 rdata7[16]
port 281 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 rdata7[17]
port 282 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 rdata7[18]
port 283 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 rdata7[19]
port 284 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 rdata7[1]
port 285 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 rdata7[20]
port 286 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 rdata7[21]
port 287 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 rdata7[22]
port 288 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 rdata7[23]
port 289 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 rdata7[24]
port 290 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 rdata7[25]
port 291 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 rdata7[26]
port 292 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 rdata7[27]
port 293 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 rdata7[28]
port 294 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 rdata7[29]
port 295 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 rdata7[2]
port 296 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 rdata7[30]
port 297 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 rdata7[31]
port 298 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 rdata7[3]
port 299 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 rdata7[4]
port 300 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 rdata7[5]
port 301 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 rdata7[6]
port 302 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 rdata7[7]
port 303 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 rdata7[8]
port 304 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 rdata7[9]
port 305 nsew signal output
rlabel metal4 s 4208 2128 4528 161616 6 vccd1
port 306 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 161616 6 vccd1
port 306 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 161616 6 vccd1
port 306 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 161616 6 vccd1
port 306 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 161616 6 vssd1
port 307 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 161616 6 vssd1
port 307 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 161616 6 vssd1
port 307 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 161616 6 vssd1
port 307 nsew ground bidirectional
rlabel metal3 s 0 3816 800 3936 6 waddr0[0]
port 308 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 waddr0[1]
port 309 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 waddr0[2]
port 310 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 waddr0[3]
port 311 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 waddr0[4]
port 312 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 waddr0[5]
port 313 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 waddr1[0]
port 314 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 waddr1[1]
port 315 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 waddr1[2]
port 316 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 waddr1[3]
port 317 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 waddr1[4]
port 318 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 waddr1[5]
port 319 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 waddr2[0]
port 320 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 waddr2[1]
port 321 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 waddr2[2]
port 322 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 waddr2[3]
port 323 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 waddr2[4]
port 324 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 waddr2[5]
port 325 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 waddr3[0]
port 326 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 waddr3[1]
port 327 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 waddr3[2]
port 328 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 waddr3[3]
port 329 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 waddr3[4]
port 330 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 waddr3[5]
port 331 nsew signal input
rlabel metal2 s 478 163200 534 164000 6 wdata0[0]
port 332 nsew signal input
rlabel metal2 s 37278 163200 37334 164000 6 wdata0[10]
port 333 nsew signal input
rlabel metal2 s 40958 163200 41014 164000 6 wdata0[11]
port 334 nsew signal input
rlabel metal2 s 44638 163200 44694 164000 6 wdata0[12]
port 335 nsew signal input
rlabel metal2 s 48318 163200 48374 164000 6 wdata0[13]
port 336 nsew signal input
rlabel metal2 s 51998 163200 52054 164000 6 wdata0[14]
port 337 nsew signal input
rlabel metal2 s 55678 163200 55734 164000 6 wdata0[15]
port 338 nsew signal input
rlabel metal2 s 59358 163200 59414 164000 6 wdata0[16]
port 339 nsew signal input
rlabel metal2 s 63038 163200 63094 164000 6 wdata0[17]
port 340 nsew signal input
rlabel metal2 s 66718 163200 66774 164000 6 wdata0[18]
port 341 nsew signal input
rlabel metal2 s 70398 163200 70454 164000 6 wdata0[19]
port 342 nsew signal input
rlabel metal2 s 4158 163200 4214 164000 6 wdata0[1]
port 343 nsew signal input
rlabel metal2 s 74078 163200 74134 164000 6 wdata0[20]
port 344 nsew signal input
rlabel metal2 s 77758 163200 77814 164000 6 wdata0[21]
port 345 nsew signal input
rlabel metal2 s 81438 163200 81494 164000 6 wdata0[22]
port 346 nsew signal input
rlabel metal2 s 85118 163200 85174 164000 6 wdata0[23]
port 347 nsew signal input
rlabel metal2 s 88798 163200 88854 164000 6 wdata0[24]
port 348 nsew signal input
rlabel metal2 s 92478 163200 92534 164000 6 wdata0[25]
port 349 nsew signal input
rlabel metal2 s 96158 163200 96214 164000 6 wdata0[26]
port 350 nsew signal input
rlabel metal2 s 99838 163200 99894 164000 6 wdata0[27]
port 351 nsew signal input
rlabel metal2 s 103518 163200 103574 164000 6 wdata0[28]
port 352 nsew signal input
rlabel metal2 s 107198 163200 107254 164000 6 wdata0[29]
port 353 nsew signal input
rlabel metal2 s 7838 163200 7894 164000 6 wdata0[2]
port 354 nsew signal input
rlabel metal2 s 110878 163200 110934 164000 6 wdata0[30]
port 355 nsew signal input
rlabel metal2 s 114558 163200 114614 164000 6 wdata0[31]
port 356 nsew signal input
rlabel metal2 s 11518 163200 11574 164000 6 wdata0[3]
port 357 nsew signal input
rlabel metal2 s 15198 163200 15254 164000 6 wdata0[4]
port 358 nsew signal input
rlabel metal2 s 18878 163200 18934 164000 6 wdata0[5]
port 359 nsew signal input
rlabel metal2 s 22558 163200 22614 164000 6 wdata0[6]
port 360 nsew signal input
rlabel metal2 s 26238 163200 26294 164000 6 wdata0[7]
port 361 nsew signal input
rlabel metal2 s 29918 163200 29974 164000 6 wdata0[8]
port 362 nsew signal input
rlabel metal2 s 33598 163200 33654 164000 6 wdata0[9]
port 363 nsew signal input
rlabel metal2 s 1398 163200 1454 164000 6 wdata1[0]
port 364 nsew signal input
rlabel metal2 s 38198 163200 38254 164000 6 wdata1[10]
port 365 nsew signal input
rlabel metal2 s 41878 163200 41934 164000 6 wdata1[11]
port 366 nsew signal input
rlabel metal2 s 45558 163200 45614 164000 6 wdata1[12]
port 367 nsew signal input
rlabel metal2 s 49238 163200 49294 164000 6 wdata1[13]
port 368 nsew signal input
rlabel metal2 s 52918 163200 52974 164000 6 wdata1[14]
port 369 nsew signal input
rlabel metal2 s 56598 163200 56654 164000 6 wdata1[15]
port 370 nsew signal input
rlabel metal2 s 60278 163200 60334 164000 6 wdata1[16]
port 371 nsew signal input
rlabel metal2 s 63958 163200 64014 164000 6 wdata1[17]
port 372 nsew signal input
rlabel metal2 s 67638 163200 67694 164000 6 wdata1[18]
port 373 nsew signal input
rlabel metal2 s 71318 163200 71374 164000 6 wdata1[19]
port 374 nsew signal input
rlabel metal2 s 5078 163200 5134 164000 6 wdata1[1]
port 375 nsew signal input
rlabel metal2 s 74998 163200 75054 164000 6 wdata1[20]
port 376 nsew signal input
rlabel metal2 s 78678 163200 78734 164000 6 wdata1[21]
port 377 nsew signal input
rlabel metal2 s 82358 163200 82414 164000 6 wdata1[22]
port 378 nsew signal input
rlabel metal2 s 86038 163200 86094 164000 6 wdata1[23]
port 379 nsew signal input
rlabel metal2 s 89718 163200 89774 164000 6 wdata1[24]
port 380 nsew signal input
rlabel metal2 s 93398 163200 93454 164000 6 wdata1[25]
port 381 nsew signal input
rlabel metal2 s 97078 163200 97134 164000 6 wdata1[26]
port 382 nsew signal input
rlabel metal2 s 100758 163200 100814 164000 6 wdata1[27]
port 383 nsew signal input
rlabel metal2 s 104438 163200 104494 164000 6 wdata1[28]
port 384 nsew signal input
rlabel metal2 s 108118 163200 108174 164000 6 wdata1[29]
port 385 nsew signal input
rlabel metal2 s 8758 163200 8814 164000 6 wdata1[2]
port 386 nsew signal input
rlabel metal2 s 111798 163200 111854 164000 6 wdata1[30]
port 387 nsew signal input
rlabel metal2 s 115478 163200 115534 164000 6 wdata1[31]
port 388 nsew signal input
rlabel metal2 s 12438 163200 12494 164000 6 wdata1[3]
port 389 nsew signal input
rlabel metal2 s 16118 163200 16174 164000 6 wdata1[4]
port 390 nsew signal input
rlabel metal2 s 19798 163200 19854 164000 6 wdata1[5]
port 391 nsew signal input
rlabel metal2 s 23478 163200 23534 164000 6 wdata1[6]
port 392 nsew signal input
rlabel metal2 s 27158 163200 27214 164000 6 wdata1[7]
port 393 nsew signal input
rlabel metal2 s 30838 163200 30894 164000 6 wdata1[8]
port 394 nsew signal input
rlabel metal2 s 34518 163200 34574 164000 6 wdata1[9]
port 395 nsew signal input
rlabel metal2 s 2318 163200 2374 164000 6 wdata2[0]
port 396 nsew signal input
rlabel metal2 s 39118 163200 39174 164000 6 wdata2[10]
port 397 nsew signal input
rlabel metal2 s 42798 163200 42854 164000 6 wdata2[11]
port 398 nsew signal input
rlabel metal2 s 46478 163200 46534 164000 6 wdata2[12]
port 399 nsew signal input
rlabel metal2 s 50158 163200 50214 164000 6 wdata2[13]
port 400 nsew signal input
rlabel metal2 s 53838 163200 53894 164000 6 wdata2[14]
port 401 nsew signal input
rlabel metal2 s 57518 163200 57574 164000 6 wdata2[15]
port 402 nsew signal input
rlabel metal2 s 61198 163200 61254 164000 6 wdata2[16]
port 403 nsew signal input
rlabel metal2 s 64878 163200 64934 164000 6 wdata2[17]
port 404 nsew signal input
rlabel metal2 s 68558 163200 68614 164000 6 wdata2[18]
port 405 nsew signal input
rlabel metal2 s 72238 163200 72294 164000 6 wdata2[19]
port 406 nsew signal input
rlabel metal2 s 5998 163200 6054 164000 6 wdata2[1]
port 407 nsew signal input
rlabel metal2 s 75918 163200 75974 164000 6 wdata2[20]
port 408 nsew signal input
rlabel metal2 s 79598 163200 79654 164000 6 wdata2[21]
port 409 nsew signal input
rlabel metal2 s 83278 163200 83334 164000 6 wdata2[22]
port 410 nsew signal input
rlabel metal2 s 86958 163200 87014 164000 6 wdata2[23]
port 411 nsew signal input
rlabel metal2 s 90638 163200 90694 164000 6 wdata2[24]
port 412 nsew signal input
rlabel metal2 s 94318 163200 94374 164000 6 wdata2[25]
port 413 nsew signal input
rlabel metal2 s 97998 163200 98054 164000 6 wdata2[26]
port 414 nsew signal input
rlabel metal2 s 101678 163200 101734 164000 6 wdata2[27]
port 415 nsew signal input
rlabel metal2 s 105358 163200 105414 164000 6 wdata2[28]
port 416 nsew signal input
rlabel metal2 s 109038 163200 109094 164000 6 wdata2[29]
port 417 nsew signal input
rlabel metal2 s 9678 163200 9734 164000 6 wdata2[2]
port 418 nsew signal input
rlabel metal2 s 112718 163200 112774 164000 6 wdata2[30]
port 419 nsew signal input
rlabel metal2 s 116398 163200 116454 164000 6 wdata2[31]
port 420 nsew signal input
rlabel metal2 s 13358 163200 13414 164000 6 wdata2[3]
port 421 nsew signal input
rlabel metal2 s 17038 163200 17094 164000 6 wdata2[4]
port 422 nsew signal input
rlabel metal2 s 20718 163200 20774 164000 6 wdata2[5]
port 423 nsew signal input
rlabel metal2 s 24398 163200 24454 164000 6 wdata2[6]
port 424 nsew signal input
rlabel metal2 s 28078 163200 28134 164000 6 wdata2[7]
port 425 nsew signal input
rlabel metal2 s 31758 163200 31814 164000 6 wdata2[8]
port 426 nsew signal input
rlabel metal2 s 35438 163200 35494 164000 6 wdata2[9]
port 427 nsew signal input
rlabel metal2 s 3238 163200 3294 164000 6 wdata3[0]
port 428 nsew signal input
rlabel metal2 s 40038 163200 40094 164000 6 wdata3[10]
port 429 nsew signal input
rlabel metal2 s 43718 163200 43774 164000 6 wdata3[11]
port 430 nsew signal input
rlabel metal2 s 47398 163200 47454 164000 6 wdata3[12]
port 431 nsew signal input
rlabel metal2 s 51078 163200 51134 164000 6 wdata3[13]
port 432 nsew signal input
rlabel metal2 s 54758 163200 54814 164000 6 wdata3[14]
port 433 nsew signal input
rlabel metal2 s 58438 163200 58494 164000 6 wdata3[15]
port 434 nsew signal input
rlabel metal2 s 62118 163200 62174 164000 6 wdata3[16]
port 435 nsew signal input
rlabel metal2 s 65798 163200 65854 164000 6 wdata3[17]
port 436 nsew signal input
rlabel metal2 s 69478 163200 69534 164000 6 wdata3[18]
port 437 nsew signal input
rlabel metal2 s 73158 163200 73214 164000 6 wdata3[19]
port 438 nsew signal input
rlabel metal2 s 6918 163200 6974 164000 6 wdata3[1]
port 439 nsew signal input
rlabel metal2 s 76838 163200 76894 164000 6 wdata3[20]
port 440 nsew signal input
rlabel metal2 s 80518 163200 80574 164000 6 wdata3[21]
port 441 nsew signal input
rlabel metal2 s 84198 163200 84254 164000 6 wdata3[22]
port 442 nsew signal input
rlabel metal2 s 87878 163200 87934 164000 6 wdata3[23]
port 443 nsew signal input
rlabel metal2 s 91558 163200 91614 164000 6 wdata3[24]
port 444 nsew signal input
rlabel metal2 s 95238 163200 95294 164000 6 wdata3[25]
port 445 nsew signal input
rlabel metal2 s 98918 163200 98974 164000 6 wdata3[26]
port 446 nsew signal input
rlabel metal2 s 102598 163200 102654 164000 6 wdata3[27]
port 447 nsew signal input
rlabel metal2 s 106278 163200 106334 164000 6 wdata3[28]
port 448 nsew signal input
rlabel metal2 s 109958 163200 110014 164000 6 wdata3[29]
port 449 nsew signal input
rlabel metal2 s 10598 163200 10654 164000 6 wdata3[2]
port 450 nsew signal input
rlabel metal2 s 113638 163200 113694 164000 6 wdata3[30]
port 451 nsew signal input
rlabel metal2 s 117318 163200 117374 164000 6 wdata3[31]
port 452 nsew signal input
rlabel metal2 s 14278 163200 14334 164000 6 wdata3[3]
port 453 nsew signal input
rlabel metal2 s 17958 163200 18014 164000 6 wdata3[4]
port 454 nsew signal input
rlabel metal2 s 21638 163200 21694 164000 6 wdata3[5]
port 455 nsew signal input
rlabel metal2 s 25318 163200 25374 164000 6 wdata3[6]
port 456 nsew signal input
rlabel metal2 s 28998 163200 29054 164000 6 wdata3[7]
port 457 nsew signal input
rlabel metal2 s 32678 163200 32734 164000 6 wdata3[8]
port 458 nsew signal input
rlabel metal2 s 36358 163200 36414 164000 6 wdata3[9]
port 459 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 wen0
port 460 nsew signal input
rlabel metal3 s 0 143216 800 143336 6 wen1
port 461 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 wen2
port 462 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 wen3
port 463 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 118000 164000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 68788904
string GDS_FILE /home/m/Builds/CaravelSoomRV-8/openlane/rf/runs/RUN_2022.11.22_22.09.39/results/signoff/RF.magic.gds
string GDS_START 182676
<< end >>

